 // connection = 0 OP mask = 15 total level = 0
cfg[0] = { 8'h2, 8'h0 }; // Enable EG test mode
cfg[1] = { 8'h20, 8'h20 }; // fill value
cfg[2] = { 8'h21, 8'h21 }; // fill value
cfg[3] = { 8'h22, 8'h22 }; // fill value
cfg[4] = { 8'h23, 8'h23 }; // fill value
cfg[5] = { 8'h24, 8'h24 }; // fill value
cfg[6] = { 8'h25, 8'h25 }; // fill value
cfg[7] = { 8'h26, 8'h26 }; // fill value
cfg[8] = { 8'h27, 8'h27 }; // fill value
cfg[9] = { 8'h28, 8'h28 }; // fill value
cfg[10] = { 8'h29, 8'h29 }; // fill value
cfg[11] = { 8'h2a, 8'h2a }; // fill value
cfg[12] = { 8'h2b, 8'h2b }; // fill value
cfg[13] = { 8'h2c, 8'h2c }; // fill value
cfg[14] = { 8'h2d, 8'h2d }; // fill value
cfg[15] = { 8'h2e, 8'h2e }; // fill value
cfg[16] = { 8'h2f, 8'h2f }; // fill value
cfg[17] = { 8'h30, 8'h30 }; // fill value
cfg[18] = { 8'h31, 8'h31 }; // fill value
cfg[19] = { 8'h32, 8'h32 }; // fill value
cfg[20] = { 8'h33, 8'h33 }; // fill value
cfg[21] = { 8'h34, 8'h34 }; // fill value
cfg[22] = { 8'h35, 8'h35 }; // fill value
cfg[23] = { 8'h36, 8'h36 }; // fill value
cfg[24] = { 8'h37, 8'h37 }; // fill value
cfg[25] = { 8'h38, 8'h38 }; // fill value
cfg[26] = { 8'h39, 8'h39 }; // fill value
cfg[27] = { 8'h3a, 8'h3a }; // fill value
cfg[28] = { 8'h3b, 8'h3b }; // fill value
cfg[29] = { 8'h3c, 8'h3c }; // fill value
cfg[30] = { 8'h3d, 8'h3d }; // fill value
cfg[31] = { 8'h3e, 8'h3e }; // fill value
cfg[32] = { 8'h3f, 8'h3f }; // fill value
cfg[33] = { 8'h80, 8'h80 }; // fill value
cfg[34] = { 8'h81, 8'h81 }; // fill value
cfg[35] = { 8'h82, 8'h82 }; // fill value
cfg[36] = { 8'h83, 8'h83 }; // fill value
cfg[37] = { 8'h84, 8'h84 }; // fill value
cfg[38] = { 8'h85, 8'h85 }; // fill value
cfg[39] = { 8'h86, 8'h86 }; // fill value
cfg[40] = { 8'h87, 8'h87 }; // fill value
cfg[41] = { 8'h88, 8'h88 }; // fill value
cfg[42] = { 8'h89, 8'h89 }; // fill value
cfg[43] = { 8'h8a, 8'h8a }; // fill value
cfg[44] = { 8'h8b, 8'h8b }; // fill value
cfg[45] = { 8'h8c, 8'h8c }; // fill value
cfg[46] = { 8'h8d, 8'h8d }; // fill value
cfg[47] = { 8'h8e, 8'h8e }; // fill value
cfg[48] = { 8'h8f, 8'h8f }; // fill value
cfg[49] = { 8'h90, 8'h90 }; // fill value
cfg[50] = { 8'h91, 8'h91 }; // fill value
cfg[51] = { 8'h92, 8'h92 }; // fill value
cfg[52] = { 8'h93, 8'h93 }; // fill value
cfg[53] = { 8'h94, 8'h94 }; // fill value
cfg[54] = { 8'h95, 8'h95 }; // fill value
cfg[55] = { 8'h96, 8'h96 }; // fill value
cfg[56] = { 8'h97, 8'h97 }; // fill value
cfg[57] = { 8'h98, 8'h98 }; // fill value
cfg[58] = { 8'h99, 8'h99 }; // fill value
cfg[59] = { 8'h9a, 8'h9a }; // fill value
cfg[60] = { 8'h9b, 8'h9b }; // fill value
cfg[61] = { 8'h9c, 8'h9c }; // fill value
cfg[62] = { 8'h9d, 8'h9d }; // fill value
cfg[63] = { 8'h9e, 8'h9e }; // fill value
cfg[64] = { 8'h9f, 8'h9f }; // fill value
cfg[65] = { 8'h28, 8'h19 }; // Key code
cfg[66] = { 8'h30, 8'he4 }; // KF
cfg[67] = { 8'h80, 8'h1f }; // Attack rate
cfg[68] = { 8'he0, 8'hf }; // Release rate
cfg[69] = { 8'h81, 8'h1f }; // Attack rate
cfg[70] = { 8'he1, 8'hf }; // Release rate
cfg[71] = { 8'h82, 8'h1f }; // Attack rate
cfg[72] = { 8'he2, 8'hf }; // Release rate
cfg[73] = { 8'h83, 8'h1f }; // Attack rate
cfg[74] = { 8'he3, 8'hf }; // Release rate
cfg[75] = { 8'h84, 8'h1f }; // Attack rate
cfg[76] = { 8'he4, 8'hf }; // Release rate
cfg[77] = { 8'h85, 8'h1f }; // Attack rate
cfg[78] = { 8'he5, 8'hf }; // Release rate
cfg[79] = { 8'h86, 8'h1f }; // Attack rate
cfg[80] = { 8'he6, 8'hf }; // Release rate
cfg[81] = { 8'h87, 8'h1f }; // Attack rate
cfg[82] = { 8'he7, 8'hf }; // Release rate
cfg[83] = { 8'h88, 8'h1f }; // Attack rate
cfg[84] = { 8'he8, 8'hf }; // Release rate
cfg[85] = { 8'h89, 8'h1f }; // Attack rate
cfg[86] = { 8'he9, 8'hf }; // Release rate
cfg[87] = { 8'h8a, 8'h1f }; // Attack rate
cfg[88] = { 8'hea, 8'hf }; // Release rate
cfg[89] = { 8'h8b, 8'h1f }; // Attack rate
cfg[90] = { 8'heb, 8'hf }; // Release rate
cfg[91] = { 8'h8c, 8'h1f }; // Attack rate
cfg[92] = { 8'hec, 8'hf }; // Release rate
cfg[93] = { 8'h8d, 8'h1f }; // Attack rate
cfg[94] = { 8'hed, 8'hf }; // Release rate
cfg[95] = { 8'h8e, 8'h1f }; // Attack rate
cfg[96] = { 8'hee, 8'hf }; // Release rate
cfg[97] = { 8'h8f, 8'h1f }; // Attack rate
cfg[98] = { 8'hef, 8'hf }; // Release rate
cfg[99] = { 8'h90, 8'h1f }; // Attack rate
cfg[100] = { 8'hf0, 8'hf }; // Release rate
cfg[101] = { 8'h91, 8'h1f }; // Attack rate
cfg[102] = { 8'hf1, 8'hf }; // Release rate
cfg[103] = { 8'h92, 8'h1f }; // Attack rate
cfg[104] = { 8'hf2, 8'hf }; // Release rate
cfg[105] = { 8'h93, 8'h1f }; // Attack rate
cfg[106] = { 8'hf3, 8'hf }; // Release rate
cfg[107] = { 8'h94, 8'h1f }; // Attack rate
cfg[108] = { 8'hf4, 8'hf }; // Release rate
cfg[109] = { 8'h95, 8'h1f }; // Attack rate
cfg[110] = { 8'hf5, 8'hf }; // Release rate
cfg[111] = { 8'h96, 8'h1f }; // Attack rate
cfg[112] = { 8'hf6, 8'hf }; // Release rate
cfg[113] = { 8'h97, 8'h1f }; // Attack rate
cfg[114] = { 8'hf7, 8'hf }; // Release rate
cfg[115] = { 8'h98, 8'h1f }; // Attack rate
cfg[116] = { 8'hf8, 8'hf }; // Release rate
cfg[117] = { 8'h99, 8'h1f }; // Attack rate
cfg[118] = { 8'hf9, 8'hf }; // Release rate
cfg[119] = { 8'h9a, 8'h1f }; // Attack rate
cfg[120] = { 8'hfa, 8'hf }; // Release rate
cfg[121] = { 8'h9b, 8'h1f }; // Attack rate
cfg[122] = { 8'hfb, 8'hf }; // Release rate
cfg[123] = { 8'h9c, 8'h1f }; // Attack rate
cfg[124] = { 8'hfc, 8'hf }; // Release rate
cfg[125] = { 8'h9d, 8'h1f }; // Attack rate
cfg[126] = { 8'hfd, 8'hf }; // Release rate
cfg[127] = { 8'h9e, 8'h1f }; // Attack rate
cfg[128] = { 8'hfe, 8'hf }; // Release rate
cfg[129] = { 8'h9f, 8'h1f }; // Attack rate
cfg[130] = { 8'hff, 8'hf }; // Release rate
cfg[131] = { 8'h8, 8'h0 }; // key off
cfg[132] = { 8'h8, 8'h1 }; // key off
cfg[133] = { 8'h8, 8'h2 }; // key off
cfg[134] = { 8'h8, 8'h3 }; // key off
cfg[135] = { 8'h8, 8'h4 }; // key off
cfg[136] = { 8'h8, 8'h5 }; // key off
cfg[137] = { 8'h8, 8'h6 }; // key off
cfg[138] = { 8'h8, 8'h7 }; // key off
cfg[139] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[140] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[141] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[142] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[143] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[144] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[145] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[146] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[147] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[148] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[149] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[150] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[151] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[152] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[153] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[154] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[155] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[156] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[157] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[158] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[159] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[160] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[161] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[162] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[163] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[164] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[165] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[166] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[167] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[168] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[169] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[170] = { 8'h1, 8'h1 }; // Gives time so keyoff works
cfg[171] = { 8'h40, 8'h1 }; // MUL
cfg[172] = { 8'h60, 8'h0 }; // TL
cfg[173] = { 8'hc0, 8'h0 }; // DT2
cfg[174] = { 8'h48, 8'h1 }; // MUL
cfg[175] = { 8'h68, 8'h0 }; // TL
cfg[176] = { 8'hc8, 8'h0 }; // DT2
cfg[177] = { 8'h50, 8'h1 }; // MUL
cfg[178] = { 8'h70, 8'h0 }; // TL
cfg[179] = { 8'hd0, 8'h0 }; // DT2
cfg[180] = { 8'h58, 8'h1 }; // MUL
cfg[181] = { 8'h78, 8'h0 }; // TL
cfg[182] = { 8'hd8, 8'h0 }; // DT2
cfg[183] = { 8'h20, 8'hc0 }; // connection
cfg[184] = { 8'h8, 8'h78 }; // key on
cfg[185] = { 8'h0, 8'h0 }; // END
