/*  This file is part of JT51.

    JT51 is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JT51 is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JT51.  If not, see <http://www.gnu.org/licenses/>.
	
	Author: Jose Tejada Gomez. Twitter: @topapate
	Version: 1.0
	Date: 27-10-2016
	*/

8'd0: pow_val <= 13'd8168;
8'd1: pow_val <= 13'd8148;
8'd2: pow_val <= 13'd8124;
8'd3: pow_val <= 13'd8104;
8'd4: pow_val <= 13'd8080;
8'd5: pow_val <= 13'd8060;
8'd6: pow_val <= 13'd8040;
8'd7: pow_val <= 13'd8016;
8'd8: pow_val <= 13'd7996;
8'd9: pow_val <= 13'd7972;
8'd10: pow_val <= 13'd7952;
8'd11: pow_val <= 13'd7932;
8'd12: pow_val <= 13'd7908;
8'd13: pow_val <= 13'd7888;
8'd14: pow_val <= 13'd7864;
8'd15: pow_val <= 13'd7844;
8'd16: pow_val <= 13'd7824;
8'd17: pow_val <= 13'd7804;
8'd18: pow_val <= 13'd7780;
8'd19: pow_val <= 13'd7760;
8'd20: pow_val <= 13'd7740;
8'd21: pow_val <= 13'd7720;
8'd22: pow_val <= 13'd7696;
8'd23: pow_val <= 13'd7676;
8'd24: pow_val <= 13'd7656;
8'd25: pow_val <= 13'd7636;
8'd26: pow_val <= 13'd7616;
8'd27: pow_val <= 13'd7592;
8'd28: pow_val <= 13'd7572;
8'd29: pow_val <= 13'd7552;
8'd30: pow_val <= 13'd7532;
8'd31: pow_val <= 13'd7512;
8'd32: pow_val <= 13'd7492;
8'd33: pow_val <= 13'd7472;
8'd34: pow_val <= 13'd7452;
8'd35: pow_val <= 13'd7432;
8'd36: pow_val <= 13'd7412;
8'd37: pow_val <= 13'd7392;
8'd38: pow_val <= 13'd7372;
8'd39: pow_val <= 13'd7352;
8'd40: pow_val <= 13'd7332;
8'd41: pow_val <= 13'd7312;
8'd42: pow_val <= 13'd7292;
8'd43: pow_val <= 13'd7272;
8'd44: pow_val <= 13'd7252;
8'd45: pow_val <= 13'd7232;
8'd46: pow_val <= 13'd7212;
8'd47: pow_val <= 13'd7192;
8'd48: pow_val <= 13'd7176;
8'd49: pow_val <= 13'd7156;
8'd50: pow_val <= 13'd7136;
8'd51: pow_val <= 13'd7116;
8'd52: pow_val <= 13'd7096;
8'd53: pow_val <= 13'd7076;
8'd54: pow_val <= 13'd7060;
8'd55: pow_val <= 13'd7040;
8'd56: pow_val <= 13'd7020;
8'd57: pow_val <= 13'd7000;
8'd58: pow_val <= 13'd6984;
8'd59: pow_val <= 13'd6964;
8'd60: pow_val <= 13'd6944;
8'd61: pow_val <= 13'd6928;
8'd62: pow_val <= 13'd6908;
8'd63: pow_val <= 13'd6888;
8'd64: pow_val <= 13'd6868;
8'd65: pow_val <= 13'd6852;
8'd66: pow_val <= 13'd6832;
8'd67: pow_val <= 13'd6816;
8'd68: pow_val <= 13'd6796;
8'd69: pow_val <= 13'd6776;
8'd70: pow_val <= 13'd6760;
8'd71: pow_val <= 13'd6740;
8'd72: pow_val <= 13'd6724;
8'd73: pow_val <= 13'd6704;
8'd74: pow_val <= 13'd6688;
8'd75: pow_val <= 13'd6668;
8'd76: pow_val <= 13'd6652;
8'd77: pow_val <= 13'd6632;
8'd78: pow_val <= 13'd6616;
8'd79: pow_val <= 13'd6596;
8'd80: pow_val <= 13'd6580;
8'd81: pow_val <= 13'd6560;
8'd82: pow_val <= 13'd6544;
8'd83: pow_val <= 13'd6524;
8'd84: pow_val <= 13'd6508;
8'd85: pow_val <= 13'd6492;
8'd86: pow_val <= 13'd6472;
8'd87: pow_val <= 13'd6456;
8'd88: pow_val <= 13'd6436;
8'd89: pow_val <= 13'd6420;
8'd90: pow_val <= 13'd6404;
8'd91: pow_val <= 13'd6384;
8'd92: pow_val <= 13'd6368;
8'd93: pow_val <= 13'd6352;
8'd94: pow_val <= 13'd6336;
8'd95: pow_val <= 13'd6316;
8'd96: pow_val <= 13'd6300;
8'd97: pow_val <= 13'd6284;
8'd98: pow_val <= 13'd6264;
8'd99: pow_val <= 13'd6248;
8'd100: pow_val <= 13'd6232;
8'd101: pow_val <= 13'd6216;
8'd102: pow_val <= 13'd6200;
8'd103: pow_val <= 13'd6180;
8'd104: pow_val <= 13'd6164;
8'd105: pow_val <= 13'd6148;
8'd106: pow_val <= 13'd6132;
8'd107: pow_val <= 13'd6116;
8'd108: pow_val <= 13'd6100;
8'd109: pow_val <= 13'd6080;
8'd110: pow_val <= 13'd6064;
8'd111: pow_val <= 13'd6048;
8'd112: pow_val <= 13'd6032;
8'd113: pow_val <= 13'd6016;
8'd114: pow_val <= 13'd6000;
8'd115: pow_val <= 13'd5984;
8'd116: pow_val <= 13'd5968;
8'd117: pow_val <= 13'd5952;
8'd118: pow_val <= 13'd5936;
8'd119: pow_val <= 13'd5920;
8'd120: pow_val <= 13'd5904;
8'd121: pow_val <= 13'd5888;
8'd122: pow_val <= 13'd5872;
8'd123: pow_val <= 13'd5856;
8'd124: pow_val <= 13'd5840;
8'd125: pow_val <= 13'd5824;
8'd126: pow_val <= 13'd5808;
8'd127: pow_val <= 13'd5792;
8'd128: pow_val <= 13'd5776;
8'd129: pow_val <= 13'd5760;
8'd130: pow_val <= 13'd5744;
8'd131: pow_val <= 13'd5732;
8'd132: pow_val <= 13'd5716;
8'd133: pow_val <= 13'd5700;
8'd134: pow_val <= 13'd5684;
8'd135: pow_val <= 13'd5668;
8'd136: pow_val <= 13'd5652;
8'd137: pow_val <= 13'd5636;
8'd138: pow_val <= 13'd5624;
8'd139: pow_val <= 13'd5608;
8'd140: pow_val <= 13'd5592;
8'd141: pow_val <= 13'd5576;
8'd142: pow_val <= 13'd5564;
8'd143: pow_val <= 13'd5548;
8'd144: pow_val <= 13'd5532;
8'd145: pow_val <= 13'd5516;
8'd146: pow_val <= 13'd5504;
8'd147: pow_val <= 13'd5488;
8'd148: pow_val <= 13'd5472;
8'd149: pow_val <= 13'd5456;
8'd150: pow_val <= 13'd5444;
8'd151: pow_val <= 13'd5428;
8'd152: pow_val <= 13'd5412;
8'd153: pow_val <= 13'd5400;
8'd154: pow_val <= 13'd5384;
8'd155: pow_val <= 13'd5368;
8'd156: pow_val <= 13'd5356;
8'd157: pow_val <= 13'd5340;
8'd158: pow_val <= 13'd5328;
8'd159: pow_val <= 13'd5312;
8'd160: pow_val <= 13'd5296;
8'd161: pow_val <= 13'd5284;
8'd162: pow_val <= 13'd5268;
8'd163: pow_val <= 13'd5256;
8'd164: pow_val <= 13'd5240;
8'd165: pow_val <= 13'd5228;
8'd166: pow_val <= 13'd5212;
8'd167: pow_val <= 13'd5200;
8'd168: pow_val <= 13'd5184;
8'd169: pow_val <= 13'd5168;
8'd170: pow_val <= 13'd5156;
8'd171: pow_val <= 13'd5144;
8'd172: pow_val <= 13'd5128;
8'd173: pow_val <= 13'd5116;
8'd174: pow_val <= 13'd5100;
8'd175: pow_val <= 13'd5088;
8'd176: pow_val <= 13'd5072;
8'd177: pow_val <= 13'd5060;
8'd178: pow_val <= 13'd5044;
8'd179: pow_val <= 13'd5032;
8'd180: pow_val <= 13'd5020;
8'd181: pow_val <= 13'd5004;
8'd182: pow_val <= 13'd4992;
8'd183: pow_val <= 13'd4976;
8'd184: pow_val <= 13'd4964;
8'd185: pow_val <= 13'd4952;
8'd186: pow_val <= 13'd4936;
8'd187: pow_val <= 13'd4924;
8'd188: pow_val <= 13'd4912;
8'd189: pow_val <= 13'd4896;
8'd190: pow_val <= 13'd4884;
8'd191: pow_val <= 13'd4872;
8'd192: pow_val <= 13'd4856;
8'd193: pow_val <= 13'd4844;
8'd194: pow_val <= 13'd4832;
8'd195: pow_val <= 13'd4820;
8'd196: pow_val <= 13'd4804;
8'd197: pow_val <= 13'd4792;
8'd198: pow_val <= 13'd4780;
8'd199: pow_val <= 13'd4768;
8'd200: pow_val <= 13'd4752;
8'd201: pow_val <= 13'd4740;
8'd202: pow_val <= 13'd4728;
8'd203: pow_val <= 13'd4716;
8'd204: pow_val <= 13'd4704;
8'd205: pow_val <= 13'd4688;
8'd206: pow_val <= 13'd4676;
8'd207: pow_val <= 13'd4664;
8'd208: pow_val <= 13'd4652;
8'd209: pow_val <= 13'd4640;
8'd210: pow_val <= 13'd4628;
8'd211: pow_val <= 13'd4616;
8'd212: pow_val <= 13'd4600;
8'd213: pow_val <= 13'd4588;
8'd214: pow_val <= 13'd4576;
8'd215: pow_val <= 13'd4564;
8'd216: pow_val <= 13'd4552;
8'd217: pow_val <= 13'd4540;
8'd218: pow_val <= 13'd4528;
8'd219: pow_val <= 13'd4516;
8'd220: pow_val <= 13'd4504;
8'd221: pow_val <= 13'd4492;
8'd222: pow_val <= 13'd4480;
8'd223: pow_val <= 13'd4468;
8'd224: pow_val <= 13'd4456;
8'd225: pow_val <= 13'd4444;
8'd226: pow_val <= 13'd4432;
8'd227: pow_val <= 13'd4420;
8'd228: pow_val <= 13'd4408;
8'd229: pow_val <= 13'd4396;
8'd230: pow_val <= 13'd4384;
8'd231: pow_val <= 13'd4372;
8'd232: pow_val <= 13'd4360;
8'd233: pow_val <= 13'd4348;
8'd234: pow_val <= 13'd4336;
8'd235: pow_val <= 13'd4324;
8'd236: pow_val <= 13'd4312;
8'd237: pow_val <= 13'd4300;
8'd238: pow_val <= 13'd4288;
8'd239: pow_val <= 13'd4276;
8'd240: pow_val <= 13'd4264;
8'd241: pow_val <= 13'd4256;
8'd242: pow_val <= 13'd4244;
8'd243: pow_val <= 13'd4232;
8'd244: pow_val <= 13'd4220;
8'd245: pow_val <= 13'd4208;
8'd246: pow_val <= 13'd4196;
8'd247: pow_val <= 13'd4184;
8'd248: pow_val <= 13'd4176;
8'd249: pow_val <= 13'd4164;
8'd250: pow_val <= 13'd4152;
8'd251: pow_val <= 13'd4140;
8'd252: pow_val <= 13'd4128;
8'd253: pow_val <= 13'd4120;
8'd254: pow_val <= 13'd4108;
8'd255: pow_val <= 13'd4096;
