 // connection = 7 OP mask = 1 total level = 0
cfg[0] = { 8'h2, 8'h0 }; // Enable EG test mode
cfg[1] = { 8'h18, 8'hff }; // LFO freq
cfg[2] = { 8'h19, 8'h7f }; // LFO AMD
cfg[3] = { 8'h19, 8'hff }; // LFO PMD
cfg[4] = { 8'h1b, 8'h1 }; // LFO waveform
cfg[5] = { 8'h28, 8'h19 }; // Key code
cfg[6] = { 8'h30, 8'he4 }; // KF
cfg[7] = { 8'he0, 8'hf }; // Release rate
cfg[8] = { 8'h60, 8'h7f }; // TL off
cfg[9] = { 8'h80, 8'h0 }; // AR as OP number
cfg[10] = { 8'he1, 8'hf }; // Release rate
cfg[11] = { 8'h61, 8'h7f }; // TL off
cfg[12] = { 8'h81, 8'h1 }; // AR as OP number
cfg[13] = { 8'he2, 8'hf }; // Release rate
cfg[14] = { 8'h62, 8'h7f }; // TL off
cfg[15] = { 8'h82, 8'h2 }; // AR as OP number
cfg[16] = { 8'he3, 8'hf }; // Release rate
cfg[17] = { 8'h63, 8'h7f }; // TL off
cfg[18] = { 8'h83, 8'h3 }; // AR as OP number
cfg[19] = { 8'he4, 8'hf }; // Release rate
cfg[20] = { 8'h64, 8'h7f }; // TL off
cfg[21] = { 8'h84, 8'h4 }; // AR as OP number
cfg[22] = { 8'he5, 8'hf }; // Release rate
cfg[23] = { 8'h65, 8'h7f }; // TL off
cfg[24] = { 8'h85, 8'h5 }; // AR as OP number
cfg[25] = { 8'he6, 8'hf }; // Release rate
cfg[26] = { 8'h66, 8'h7f }; // TL off
cfg[27] = { 8'h86, 8'h6 }; // AR as OP number
cfg[28] = { 8'he7, 8'hf }; // Release rate
cfg[29] = { 8'h67, 8'h7f }; // TL off
cfg[30] = { 8'h87, 8'h7 }; // AR as OP number
cfg[31] = { 8'he8, 8'hf }; // Release rate
cfg[32] = { 8'h68, 8'h7f }; // TL off
cfg[33] = { 8'h88, 8'h8 }; // AR as OP number
cfg[34] = { 8'he9, 8'hf }; // Release rate
cfg[35] = { 8'h69, 8'h7f }; // TL off
cfg[36] = { 8'h89, 8'h9 }; // AR as OP number
cfg[37] = { 8'hea, 8'hf }; // Release rate
cfg[38] = { 8'h6a, 8'h7f }; // TL off
cfg[39] = { 8'h8a, 8'ha }; // AR as OP number
cfg[40] = { 8'heb, 8'hf }; // Release rate
cfg[41] = { 8'h6b, 8'h7f }; // TL off
cfg[42] = { 8'h8b, 8'hb }; // AR as OP number
cfg[43] = { 8'hec, 8'hf }; // Release rate
cfg[44] = { 8'h6c, 8'h7f }; // TL off
cfg[45] = { 8'h8c, 8'hc }; // AR as OP number
cfg[46] = { 8'hed, 8'hf }; // Release rate
cfg[47] = { 8'h6d, 8'h7f }; // TL off
cfg[48] = { 8'h8d, 8'hd }; // AR as OP number
cfg[49] = { 8'hee, 8'hf }; // Release rate
cfg[50] = { 8'h6e, 8'h7f }; // TL off
cfg[51] = { 8'h8e, 8'he }; // AR as OP number
cfg[52] = { 8'hef, 8'hf }; // Release rate
cfg[53] = { 8'h6f, 8'h7f }; // TL off
cfg[54] = { 8'h8f, 8'hf }; // AR as OP number
cfg[55] = { 8'hf0, 8'hf }; // Release rate
cfg[56] = { 8'h70, 8'h7f }; // TL off
cfg[57] = { 8'h90, 8'h10 }; // AR as OP number
cfg[58] = { 8'hf1, 8'hf }; // Release rate
cfg[59] = { 8'h71, 8'h7f }; // TL off
cfg[60] = { 8'h91, 8'h11 }; // AR as OP number
cfg[61] = { 8'hf2, 8'hf }; // Release rate
cfg[62] = { 8'h72, 8'h7f }; // TL off
cfg[63] = { 8'h92, 8'h12 }; // AR as OP number
cfg[64] = { 8'hf3, 8'hf }; // Release rate
cfg[65] = { 8'h73, 8'h7f }; // TL off
cfg[66] = { 8'h93, 8'h13 }; // AR as OP number
cfg[67] = { 8'hf4, 8'hf }; // Release rate
cfg[68] = { 8'h74, 8'h7f }; // TL off
cfg[69] = { 8'h94, 8'h14 }; // AR as OP number
cfg[70] = { 8'hf5, 8'hf }; // Release rate
cfg[71] = { 8'h75, 8'h7f }; // TL off
cfg[72] = { 8'h95, 8'h15 }; // AR as OP number
cfg[73] = { 8'hf6, 8'hf }; // Release rate
cfg[74] = { 8'h76, 8'h7f }; // TL off
cfg[75] = { 8'h96, 8'h16 }; // AR as OP number
cfg[76] = { 8'hf7, 8'hf }; // Release rate
cfg[77] = { 8'h77, 8'h7f }; // TL off
cfg[78] = { 8'h97, 8'h17 }; // AR as OP number
cfg[79] = { 8'hf8, 8'hf }; // Release rate
cfg[80] = { 8'h78, 8'h7f }; // TL off
cfg[81] = { 8'h98, 8'h18 }; // AR as OP number
cfg[82] = { 8'hf9, 8'hf }; // Release rate
cfg[83] = { 8'h79, 8'h7f }; // TL off
cfg[84] = { 8'h99, 8'h19 }; // AR as OP number
cfg[85] = { 8'hfa, 8'hf }; // Release rate
cfg[86] = { 8'h7a, 8'h7f }; // TL off
cfg[87] = { 8'h9a, 8'h1a }; // AR as OP number
cfg[88] = { 8'hfb, 8'hf }; // Release rate
cfg[89] = { 8'h7b, 8'h7f }; // TL off
cfg[90] = { 8'h9b, 8'h1b }; // AR as OP number
cfg[91] = { 8'hfc, 8'hf }; // Release rate
cfg[92] = { 8'h7c, 8'h7f }; // TL off
cfg[93] = { 8'h9c, 8'h1c }; // AR as OP number
cfg[94] = { 8'hfd, 8'hf }; // Release rate
cfg[95] = { 8'h7d, 8'h7f }; // TL off
cfg[96] = { 8'h9d, 8'h1d }; // AR as OP number
cfg[97] = { 8'hfe, 8'hf }; // Release rate
cfg[98] = { 8'h7e, 8'h7f }; // TL off
cfg[99] = { 8'h9e, 8'h1e }; // AR as OP number
cfg[100] = { 8'hff, 8'hf }; // Release rate
cfg[101] = { 8'h7f, 8'h7f }; // TL off
cfg[102] = { 8'h9f, 8'h1f }; // AR as OP number
cfg[103] = { 8'h40, 8'h1 }; // MUL
cfg[104] = { 8'h60, 8'h0 }; // TL
cfg[105] = { 8'h48, 8'h1 }; // MUL
cfg[106] = { 8'h50, 8'h1 }; // MUL
cfg[107] = { 8'h58, 8'h1 }; // MUL
cfg[108] = { 8'h8, 8'h0 }; // key off
cfg[109] = { 8'h20, 8'h7 };
cfg[110] = { 8'h8, 8'h1 }; // key off
cfg[111] = { 8'h21, 8'h7 };
cfg[112] = { 8'h8, 8'h2 }; // key off
cfg[113] = { 8'h22, 8'h7 };
cfg[114] = { 8'h8, 8'h3 }; // key off
cfg[115] = { 8'h23, 8'h7 };
cfg[116] = { 8'h8, 8'h4 }; // key off
cfg[117] = { 8'h24, 8'h7 };
cfg[118] = { 8'h8, 8'h5 }; // key off
cfg[119] = { 8'h25, 8'h7 };
cfg[120] = { 8'h8, 8'h6 }; // key off
cfg[121] = { 8'h26, 8'h7 };
cfg[122] = { 8'h8, 8'h7 }; // key off
cfg[123] = { 8'h27, 8'h7 };
cfg[124] = { 8'h20, 8'hcf }; // connection
cfg[125] = { 8'h38, 8'h2 }; // PMS/AMS
cfg[126] = { 8'h80, 8'h1f }; // KS/AR
cfg[127] = { 8'ha0, 8'h80 }; // AMSEN / D1R rate
cfg[128] = { 8'hc0, 8'h0 }; // DT2 / D2R rate
cfg[129] = { 8'he0, 8'hcf }; // D1L/RR
cfg[130] = { 8'h88, 8'h1f }; // KS/AR
cfg[131] = { 8'ha8, 8'h80 }; // AMSEN / D1R rate
cfg[132] = { 8'hc8, 8'h0 }; // DT2 / D2R rate
cfg[133] = { 8'he8, 8'hcf }; // D1L/RR
cfg[134] = { 8'h90, 8'h1f }; // KS/AR
cfg[135] = { 8'hb0, 8'h80 }; // AMSEN / D1R rate
cfg[136] = { 8'hd0, 8'h0 }; // DT2 / D2R rate
cfg[137] = { 8'hf0, 8'hcf }; // D1L/RR
cfg[138] = { 8'h98, 8'h1f }; // KS/AR
cfg[139] = { 8'hb8, 8'h80 }; // AMSEN / D1R rate
cfg[140] = { 8'hd8, 8'h0 }; // DT2 / D2R rate
cfg[141] = { 8'hf8, 8'hcf }; // D1L/RR
cfg[142] = { 8'h8, 8'h8 }; // key on
cfg[143] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[144] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[145] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[146] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[147] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[148] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[149] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[150] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[151] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[152] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[153] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[154] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[155] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[156] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[157] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[158] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[159] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[160] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[161] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[162] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[163] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[164] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[165] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[166] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[167] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[168] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[169] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[170] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[171] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[172] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[173] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[174] = { 8'h1, 8'h1 }; // Gives time so sound can start
cfg[175] = { 8'h0, 8'h0 }; // END
