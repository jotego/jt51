/*  This file is part of JT51.

    JT51 is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JT51 is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JT51.  If not, see <http://www.gnu.org/licenses/>.
	
	Author: Jose Tejada Gomez. Twitter: @topapate
	Version: 1.0
	Date: 27-10-2016
	*/
	
8'd0: log_val <= 12'd2137;
8'd1: log_val <= 12'd1731;
8'd2: log_val <= 12'd1543;
8'd3: log_val <= 12'd1419;
8'd4: log_val <= 12'd1326;
8'd5: log_val <= 12'd1252;
8'd6: log_val <= 12'd1190;
8'd7: log_val <= 12'd1137;
8'd8: log_val <= 12'd1091;
8'd9: log_val <= 12'd1050;
8'd10: log_val <= 12'd1013;
8'd11: log_val <= 12'd979;
8'd12: log_val <= 12'd949;
8'd13: log_val <= 12'd920;
8'd14: log_val <= 12'd894;
8'd15: log_val <= 12'd869;
8'd16: log_val <= 12'd846;
8'd17: log_val <= 12'd825;
8'd18: log_val <= 12'd804;
8'd19: log_val <= 12'd785;
8'd20: log_val <= 12'd767;
8'd21: log_val <= 12'd749;
8'd22: log_val <= 12'd732;
8'd23: log_val <= 12'd717;
8'd24: log_val <= 12'd701;
8'd25: log_val <= 12'd687;
8'd26: log_val <= 12'd672;
8'd27: log_val <= 12'd659;
8'd28: log_val <= 12'd646;
8'd29: log_val <= 12'd633;
8'd30: log_val <= 12'd621;
8'd31: log_val <= 12'd609;
8'd32: log_val <= 12'd598;
8'd33: log_val <= 12'd587;
8'd34: log_val <= 12'd576;
8'd35: log_val <= 12'd566;
8'd36: log_val <= 12'd556;
8'd37: log_val <= 12'd546;
8'd38: log_val <= 12'd536;
8'd39: log_val <= 12'd527;
8'd40: log_val <= 12'd518;
8'd41: log_val <= 12'd509;
8'd42: log_val <= 12'd501;
8'd43: log_val <= 12'd492;
8'd44: log_val <= 12'd484;
8'd45: log_val <= 12'd476;
8'd46: log_val <= 12'd468;
8'd47: log_val <= 12'd461;
8'd48: log_val <= 12'd453;
8'd49: log_val <= 12'd446;
8'd50: log_val <= 12'd439;
8'd51: log_val <= 12'd432;
8'd52: log_val <= 12'd425;
8'd53: log_val <= 12'd418;
8'd54: log_val <= 12'd411;
8'd55: log_val <= 12'd405;
8'd56: log_val <= 12'd399;
8'd57: log_val <= 12'd392;
8'd58: log_val <= 12'd386;
8'd59: log_val <= 12'd380;
8'd60: log_val <= 12'd375;
8'd61: log_val <= 12'd369;
8'd62: log_val <= 12'd363;
8'd63: log_val <= 12'd358;
8'd64: log_val <= 12'd352;
8'd65: log_val <= 12'd347;
8'd66: log_val <= 12'd341;
8'd67: log_val <= 12'd336;
8'd68: log_val <= 12'd331;
8'd69: log_val <= 12'd326;
8'd70: log_val <= 12'd321;
8'd71: log_val <= 12'd316;
8'd72: log_val <= 12'd311;
8'd73: log_val <= 12'd307;
8'd74: log_val <= 12'd302;
8'd75: log_val <= 12'd297;
8'd76: log_val <= 12'd293;
8'd77: log_val <= 12'd289;
8'd78: log_val <= 12'd284;
8'd79: log_val <= 12'd280;
8'd80: log_val <= 12'd276;
8'd81: log_val <= 12'd271;
8'd82: log_val <= 12'd267;
8'd83: log_val <= 12'd263;
8'd84: log_val <= 12'd259;
8'd85: log_val <= 12'd255;
8'd86: log_val <= 12'd251;
8'd87: log_val <= 12'd248;
8'd88: log_val <= 12'd244;
8'd89: log_val <= 12'd240;
8'd90: log_val <= 12'd236;
8'd91: log_val <= 12'd233;
8'd92: log_val <= 12'd229;
8'd93: log_val <= 12'd226;
8'd94: log_val <= 12'd222;
8'd95: log_val <= 12'd219;
8'd96: log_val <= 12'd215;
8'd97: log_val <= 12'd212;
8'd98: log_val <= 12'd209;
8'd99: log_val <= 12'd205;
8'd100: log_val <= 12'd202;
8'd101: log_val <= 12'd199;
8'd102: log_val <= 12'd196;
8'd103: log_val <= 12'd193;
8'd104: log_val <= 12'd190;
8'd105: log_val <= 12'd187;
8'd106: log_val <= 12'd184;
8'd107: log_val <= 12'd181;
8'd108: log_val <= 12'd178;
8'd109: log_val <= 12'd175;
8'd110: log_val <= 12'd172;
8'd111: log_val <= 12'd169;
8'd112: log_val <= 12'd167;
8'd113: log_val <= 12'd164;
8'd114: log_val <= 12'd161;
8'd115: log_val <= 12'd159;
8'd116: log_val <= 12'd156;
8'd117: log_val <= 12'd153;
8'd118: log_val <= 12'd151;
8'd119: log_val <= 12'd148;
8'd120: log_val <= 12'd146;
8'd121: log_val <= 12'd143;
8'd122: log_val <= 12'd141;
8'd123: log_val <= 12'd138;
8'd124: log_val <= 12'd136;
8'd125: log_val <= 12'd134;
8'd126: log_val <= 12'd131;
8'd127: log_val <= 12'd129;
8'd128: log_val <= 12'd127;
8'd129: log_val <= 12'd125;
8'd130: log_val <= 12'd122;
8'd131: log_val <= 12'd120;
8'd132: log_val <= 12'd118;
8'd133: log_val <= 12'd116;
8'd134: log_val <= 12'd114;
8'd135: log_val <= 12'd112;
8'd136: log_val <= 12'd110;
8'd137: log_val <= 12'd108;
8'd138: log_val <= 12'd106;
8'd139: log_val <= 12'd104;
8'd140: log_val <= 12'd102;
8'd141: log_val <= 12'd100;
8'd142: log_val <= 12'd98;
8'd143: log_val <= 12'd96;
8'd144: log_val <= 12'd94;
8'd145: log_val <= 12'd92;
8'd146: log_val <= 12'd91;
8'd147: log_val <= 12'd89;
8'd148: log_val <= 12'd87;
8'd149: log_val <= 12'd85;
8'd150: log_val <= 12'd83;
8'd151: log_val <= 12'd82;
8'd152: log_val <= 12'd80;
8'd153: log_val <= 12'd78;
8'd154: log_val <= 12'd77;
8'd155: log_val <= 12'd75;
8'd156: log_val <= 12'd74;
8'd157: log_val <= 12'd72;
8'd158: log_val <= 12'd70;
8'd159: log_val <= 12'd69;
8'd160: log_val <= 12'd67;
8'd161: log_val <= 12'd66;
8'd162: log_val <= 12'd64;
8'd163: log_val <= 12'd63;
8'd164: log_val <= 12'd62;
8'd165: log_val <= 12'd60;
8'd166: log_val <= 12'd59;
8'd167: log_val <= 12'd57;
8'd168: log_val <= 12'd56;
8'd169: log_val <= 12'd55;
8'd170: log_val <= 12'd53;
8'd171: log_val <= 12'd52;
8'd172: log_val <= 12'd51;
8'd173: log_val <= 12'd49;
8'd174: log_val <= 12'd48;
8'd175: log_val <= 12'd47;
8'd176: log_val <= 12'd46;
8'd177: log_val <= 12'd45;
8'd178: log_val <= 12'd43;
8'd179: log_val <= 12'd42;
8'd180: log_val <= 12'd41;
8'd181: log_val <= 12'd40;
8'd182: log_val <= 12'd39;
8'd183: log_val <= 12'd38;
8'd184: log_val <= 12'd37;
8'd185: log_val <= 12'd36;
8'd186: log_val <= 12'd35;
8'd187: log_val <= 12'd34;
8'd188: log_val <= 12'd33;
8'd189: log_val <= 12'd32;
8'd190: log_val <= 12'd31;
8'd191: log_val <= 12'd30;
8'd192: log_val <= 12'd29;
8'd193: log_val <= 12'd28;
8'd194: log_val <= 12'd27;
8'd195: log_val <= 12'd26;
8'd196: log_val <= 12'd25;
8'd197: log_val <= 12'd24;
8'd198: log_val <= 12'd23;
8'd199: log_val <= 12'd23;
8'd200: log_val <= 12'd22;
8'd201: log_val <= 12'd21;
8'd202: log_val <= 12'd20;
8'd203: log_val <= 12'd20;
8'd204: log_val <= 12'd19;
8'd205: log_val <= 12'd18;
8'd206: log_val <= 12'd17;
8'd207: log_val <= 12'd17;
8'd208: log_val <= 12'd16;
8'd209: log_val <= 12'd15;
8'd210: log_val <= 12'd15;
8'd211: log_val <= 12'd14;
8'd212: log_val <= 12'd13;
8'd213: log_val <= 12'd13;
8'd214: log_val <= 12'd12;
8'd215: log_val <= 12'd12;
8'd216: log_val <= 12'd11;
8'd217: log_val <= 12'd10;
8'd218: log_val <= 12'd10;
8'd219: log_val <= 12'd9;
8'd220: log_val <= 12'd9;
8'd221: log_val <= 12'd8;
8'd222: log_val <= 12'd8;
8'd223: log_val <= 12'd7;
8'd224: log_val <= 12'd7;
8'd225: log_val <= 12'd7;
8'd226: log_val <= 12'd6;
8'd227: log_val <= 12'd6;
8'd228: log_val <= 12'd5;
8'd229: log_val <= 12'd5;
8'd230: log_val <= 12'd5;
8'd231: log_val <= 12'd4;
8'd232: log_val <= 12'd4;
8'd233: log_val <= 12'd4;
8'd234: log_val <= 12'd3;
8'd235: log_val <= 12'd3;
8'd236: log_val <= 12'd3;
8'd237: log_val <= 12'd2;
8'd238: log_val <= 12'd2;
8'd239: log_val <= 12'd2;
8'd240: log_val <= 12'd2;
8'd241: log_val <= 12'd1;
8'd242: log_val <= 12'd1;
8'd243: log_val <= 12'd1;
8'd244: log_val <= 12'd1;
8'd245: log_val <= 12'd1;
8'd246: log_val <= 12'd1;
8'd247: log_val <= 12'd1;
8'd248: log_val <= 12'd0;
8'd249: log_val <= 12'd0;
8'd250: log_val <= 12'd0;
8'd251: log_val <= 12'd0;
8'd252: log_val <= 12'd0;
8'd253: log_val <= 12'd0;
8'd254: log_val <= 12'd0;
8'd255: log_val <= 12'd0;
