/*  This file is part of JT51.

    JT51 is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JT51 is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JT51.  If not, see <http://www.gnu.org/licenses/>.

	Author: Jose Tejada Gomez. Twitter: @topapate
	Version: 1.0
	Date: 27-10-2016
	*/


module jt51_phinc_rom(
	// input				clk,
	input  		[9:0]	keycode,
	output reg	[11:0]	phinc
);

always @(*) begin : read_lut
	case( keycode )
        10'd0   : phinc={ 12'd1299 };
        10'd1   : phinc={ 12'd1300 };
        10'd2   : phinc={ 12'd1301 };
        10'd3   : phinc={ 12'd1302 };
        10'd4   : phinc={ 12'd1303 };
        10'd5   : phinc={ 12'd1304 };
        10'd6   : phinc={ 12'd1305 };
        10'd7   : phinc={ 12'd1306 };
        10'd8   : phinc={ 12'd1308 };
        10'd9   : phinc={ 12'd1309 };
        10'd10  : phinc={ 12'd1310 };
        10'd11  : phinc={ 12'd1311 };
        10'd12  : phinc={ 12'd1313 };
        10'd13  : phinc={ 12'd1314 };
        10'd14  : phinc={ 12'd1315 };
        10'd15  : phinc={ 12'd1316 };
        10'd16  : phinc={ 12'd1318 };
        10'd17  : phinc={ 12'd1319 };
        10'd18  : phinc={ 12'd1320 };
        10'd19  : phinc={ 12'd1321 };
        10'd20  : phinc={ 12'd1322 };
        10'd21  : phinc={ 12'd1323 };
        10'd22  : phinc={ 12'd1324 };
        10'd23  : phinc={ 12'd1325 };
        10'd24  : phinc={ 12'd1327 };
        10'd25  : phinc={ 12'd1328 };
        10'd26  : phinc={ 12'd1329 };
        10'd27  : phinc={ 12'd1330 };
        10'd28  : phinc={ 12'd1332 };
        10'd29  : phinc={ 12'd1333 };
        10'd30  : phinc={ 12'd1334 };
        10'd31  : phinc={ 12'd1335 };
        10'd32  : phinc={ 12'd1337 };
        10'd33  : phinc={ 12'd1338 };
        10'd34  : phinc={ 12'd1339 };
        10'd35  : phinc={ 12'd1340 };
        10'd36  : phinc={ 12'd1341 };
        10'd37  : phinc={ 12'd1342 };
        10'd38  : phinc={ 12'd1343 };
        10'd39  : phinc={ 12'd1344 };
        10'd40  : phinc={ 12'd1346 };
        10'd41  : phinc={ 12'd1347 };
        10'd42  : phinc={ 12'd1348 };
        10'd43  : phinc={ 12'd1349 };
        10'd44  : phinc={ 12'd1351 };
        10'd45  : phinc={ 12'd1352 };
        10'd46  : phinc={ 12'd1353 };
        10'd47  : phinc={ 12'd1354 };
        10'd48  : phinc={ 12'd1356 };
        10'd49  : phinc={ 12'd1357 };
        10'd50  : phinc={ 12'd1358 };
        10'd51  : phinc={ 12'd1359 };
        10'd52  : phinc={ 12'd1361 };
        10'd53  : phinc={ 12'd1362 };
        10'd54  : phinc={ 12'd1363 };
        10'd55  : phinc={ 12'd1364 };
        10'd56  : phinc={ 12'd1366 };
        10'd57  : phinc={ 12'd1367 };
        10'd58  : phinc={ 12'd1368 };
        10'd59  : phinc={ 12'd1369 };
        10'd60  : phinc={ 12'd1371 };
        10'd61  : phinc={ 12'd1372 };
        10'd62  : phinc={ 12'd1373 };
        10'd63  : phinc={ 12'd1374 };
        10'd64  : phinc={ 12'd1376 };
        10'd65  : phinc={ 12'd1377 };
        10'd66  : phinc={ 12'd1378 };
        10'd67  : phinc={ 12'd1379 };
        10'd68  : phinc={ 12'd1381 };
        10'd69  : phinc={ 12'd1382 };
        10'd70  : phinc={ 12'd1383 };
        10'd71  : phinc={ 12'd1384 };
        10'd72  : phinc={ 12'd1386 };
        10'd73  : phinc={ 12'd1387 };
        10'd74  : phinc={ 12'd1388 };
        10'd75  : phinc={ 12'd1389 };
        10'd76  : phinc={ 12'd1391 };
        10'd77  : phinc={ 12'd1392 };
        10'd78  : phinc={ 12'd1393 };
        10'd79  : phinc={ 12'd1394 };
        10'd80  : phinc={ 12'd1396 };
        10'd81  : phinc={ 12'd1397 };
        10'd82  : phinc={ 12'd1398 };
        10'd83  : phinc={ 12'd1399 };
        10'd84  : phinc={ 12'd1401 };
        10'd85  : phinc={ 12'd1402 };
        10'd86  : phinc={ 12'd1403 };
        10'd87  : phinc={ 12'd1404 };
        10'd88  : phinc={ 12'd1406 };
        10'd89  : phinc={ 12'd1407 };
        10'd90  : phinc={ 12'd1408 };
        10'd91  : phinc={ 12'd1409 };
        10'd92  : phinc={ 12'd1411 };
        10'd93  : phinc={ 12'd1412 };
        10'd94  : phinc={ 12'd1413 };
        10'd95  : phinc={ 12'd1414 };
        10'd96  : phinc={ 12'd1416 };
        10'd97  : phinc={ 12'd1417 };
        10'd98  : phinc={ 12'd1418 };
        10'd99  : phinc={ 12'd1419 };
        10'd100 : phinc={ 12'd1421 };
        10'd101 : phinc={ 12'd1422 };
        10'd102 : phinc={ 12'd1423 };
        10'd103 : phinc={ 12'd1424 };
        10'd104 : phinc={ 12'd1426 };
        10'd105 : phinc={ 12'd1427 };
        10'd106 : phinc={ 12'd1429 };
        10'd107 : phinc={ 12'd1430 };
        10'd108 : phinc={ 12'd1431 };
        10'd109 : phinc={ 12'd1432 };
        10'd110 : phinc={ 12'd1434 };
        10'd111 : phinc={ 12'd1435 };
        10'd112 : phinc={ 12'd1437 };
        10'd113 : phinc={ 12'd1438 };
        10'd114 : phinc={ 12'd1439 };
        10'd115 : phinc={ 12'd1440 };
        10'd116 : phinc={ 12'd1442 };
        10'd117 : phinc={ 12'd1443 };
        10'd118 : phinc={ 12'd1444 };
        10'd119 : phinc={ 12'd1445 };
        10'd120 : phinc={ 12'd1447 };
        10'd121 : phinc={ 12'd1448 };
        10'd122 : phinc={ 12'd1449 };
        10'd123 : phinc={ 12'd1450 };
        10'd124 : phinc={ 12'd1452 };
        10'd125 : phinc={ 12'd1453 };
        10'd126 : phinc={ 12'd1454 };
        10'd127 : phinc={ 12'd1455 };
        10'd128 : phinc={ 12'd1458 };
        10'd129 : phinc={ 12'd1459 };
        10'd130 : phinc={ 12'd1460 };
        10'd131 : phinc={ 12'd1461 };
        10'd132 : phinc={ 12'd1463 };
        10'd133 : phinc={ 12'd1464 };
        10'd134 : phinc={ 12'd1465 };
        10'd135 : phinc={ 12'd1466 };
        10'd136 : phinc={ 12'd1468 };
        10'd137 : phinc={ 12'd1469 };
        10'd138 : phinc={ 12'd1471 };
        10'd139 : phinc={ 12'd1472 };
        10'd140 : phinc={ 12'd1473 };
        10'd141 : phinc={ 12'd1474 };
        10'd142 : phinc={ 12'd1476 };
        10'd143 : phinc={ 12'd1477 };
        10'd144 : phinc={ 12'd1479 };
        10'd145 : phinc={ 12'd1480 };
        10'd146 : phinc={ 12'd1481 };
        10'd147 : phinc={ 12'd1482 };
        10'd148 : phinc={ 12'd1484 };
        10'd149 : phinc={ 12'd1485 };
        10'd150 : phinc={ 12'd1486 };
        10'd151 : phinc={ 12'd1487 };
        10'd152 : phinc={ 12'd1489 };
        10'd153 : phinc={ 12'd1490 };
        10'd154 : phinc={ 12'd1492 };
        10'd155 : phinc={ 12'd1493 };
        10'd156 : phinc={ 12'd1494 };
        10'd157 : phinc={ 12'd1495 };
        10'd158 : phinc={ 12'd1497 };
        10'd159 : phinc={ 12'd1498 };
        10'd160 : phinc={ 12'd1501 };
        10'd161 : phinc={ 12'd1502 };
        10'd162 : phinc={ 12'd1503 };
        10'd163 : phinc={ 12'd1504 };
        10'd164 : phinc={ 12'd1506 };
        10'd165 : phinc={ 12'd1507 };
        10'd166 : phinc={ 12'd1509 };
        10'd167 : phinc={ 12'd1510 };
        10'd168 : phinc={ 12'd1512 };
        10'd169 : phinc={ 12'd1513 };
        10'd170 : phinc={ 12'd1514 };
        10'd171 : phinc={ 12'd1515 };
        10'd172 : phinc={ 12'd1517 };
        10'd173 : phinc={ 12'd1518 };
        10'd174 : phinc={ 12'd1520 };
        10'd175 : phinc={ 12'd1521 };
        10'd176 : phinc={ 12'd1523 };
        10'd177 : phinc={ 12'd1524 };
        10'd178 : phinc={ 12'd1525 };
        10'd179 : phinc={ 12'd1526 };
        10'd180 : phinc={ 12'd1528 };
        10'd181 : phinc={ 12'd1529 };
        10'd182 : phinc={ 12'd1531 };
        10'd183 : phinc={ 12'd1532 };
        10'd184 : phinc={ 12'd1534 };
        10'd185 : phinc={ 12'd1535 };
        10'd186 : phinc={ 12'd1536 };
        10'd187 : phinc={ 12'd1537 };
        10'd188 : phinc={ 12'd1539 };
        10'd189 : phinc={ 12'd1540 };
        10'd190 : phinc={ 12'd1542 };
        10'd191 : phinc={ 12'd1543 };
        10'd192 : phinc={ 12'd0 };
        10'd193 : phinc={ 12'd2 };
        10'd194 : phinc={ 12'd4 };
        10'd195 : phinc={ 12'd6 };
        10'd196 : phinc={ 12'd4 };
        10'd197 : phinc={ 12'd6 };
        10'd198 : phinc={ 12'd8 };
        10'd199 : phinc={ 12'd10 };
        10'd200 : phinc={ 12'd9 };
        10'd201 : phinc={ 12'd11 };
        10'd202 : phinc={ 12'd13 };
        10'd203 : phinc={ 12'd15 };
        10'd204 : phinc={ 12'd15 };
        10'd205 : phinc={ 12'd17 };
        10'd206 : phinc={ 12'd19 };
        10'd207 : phinc={ 12'd21 };
        10'd208 : phinc={ 12'd0 };
        10'd209 : phinc={ 12'd2 };
        10'd210 : phinc={ 12'd4 };
        10'd211 : phinc={ 12'd6 };
        10'd212 : phinc={ 12'd4 };
        10'd213 : phinc={ 12'd6 };
        10'd214 : phinc={ 12'd8 };
        10'd215 : phinc={ 12'd10 };
        10'd216 : phinc={ 12'd9 };
        10'd217 : phinc={ 12'd11 };
        10'd218 : phinc={ 12'd13 };
        10'd219 : phinc={ 12'd15 };
        10'd220 : phinc={ 12'd15 };
        10'd221 : phinc={ 12'd17 };
        10'd222 : phinc={ 12'd19 };
        10'd223 : phinc={ 12'd21 };
        10'd224 : phinc={ 12'd0 };
        10'd225 : phinc={ 12'd2 };
        10'd226 : phinc={ 12'd4 };
        10'd227 : phinc={ 12'd6 };
        10'd228 : phinc={ 12'd4 };
        10'd229 : phinc={ 12'd6 };
        10'd230 : phinc={ 12'd8 };
        10'd231 : phinc={ 12'd10 };
        10'd232 : phinc={ 12'd9 };
        10'd233 : phinc={ 12'd11 };
        10'd234 : phinc={ 12'd13 };
        10'd235 : phinc={ 12'd15 };
        10'd236 : phinc={ 12'd15 };
        10'd237 : phinc={ 12'd17 };
        10'd238 : phinc={ 12'd19 };
        10'd239 : phinc={ 12'd21 };
        10'd240 : phinc={ 12'd0 };
        10'd241 : phinc={ 12'd2 };
        10'd242 : phinc={ 12'd4 };
        10'd243 : phinc={ 12'd6 };
        10'd244 : phinc={ 12'd4 };
        10'd245 : phinc={ 12'd6 };
        10'd246 : phinc={ 12'd8 };
        10'd247 : phinc={ 12'd10 };
        10'd248 : phinc={ 12'd9 };
        10'd249 : phinc={ 12'd11 };
        10'd250 : phinc={ 12'd13 };
        10'd251 : phinc={ 12'd15 };
        10'd252 : phinc={ 12'd15 };
        10'd253 : phinc={ 12'd17 };
        10'd254 : phinc={ 12'd19 };
        10'd255 : phinc={ 12'd21 };
        10'd256 : phinc={ 12'd1545 };
        10'd257 : phinc={ 12'd1546 };
        10'd258 : phinc={ 12'd1547 };
        10'd259 : phinc={ 12'd1548 };
        10'd260 : phinc={ 12'd1550 };
        10'd261 : phinc={ 12'd1551 };
        10'd262 : phinc={ 12'd1553 };
        10'd263 : phinc={ 12'd1554 };
        10'd264 : phinc={ 12'd1556 };
        10'd265 : phinc={ 12'd1557 };
        10'd266 : phinc={ 12'd1558 };
        10'd267 : phinc={ 12'd1559 };
        10'd268 : phinc={ 12'd1561 };
        10'd269 : phinc={ 12'd1562 };
        10'd270 : phinc={ 12'd1564 };
        10'd271 : phinc={ 12'd1565 };
        10'd272 : phinc={ 12'd1567 };
        10'd273 : phinc={ 12'd1568 };
        10'd274 : phinc={ 12'd1569 };
        10'd275 : phinc={ 12'd1570 };
        10'd276 : phinc={ 12'd1572 };
        10'd277 : phinc={ 12'd1573 };
        10'd278 : phinc={ 12'd1575 };
        10'd279 : phinc={ 12'd1576 };
        10'd280 : phinc={ 12'd1578 };
        10'd281 : phinc={ 12'd1579 };
        10'd282 : phinc={ 12'd1580 };
        10'd283 : phinc={ 12'd1581 };
        10'd284 : phinc={ 12'd1583 };
        10'd285 : phinc={ 12'd1584 };
        10'd286 : phinc={ 12'd1586 };
        10'd287 : phinc={ 12'd1587 };
        10'd288 : phinc={ 12'd1590 };
        10'd289 : phinc={ 12'd1591 };
        10'd290 : phinc={ 12'd1592 };
        10'd291 : phinc={ 12'd1593 };
        10'd292 : phinc={ 12'd1595 };
        10'd293 : phinc={ 12'd1596 };
        10'd294 : phinc={ 12'd1598 };
        10'd295 : phinc={ 12'd1599 };
        10'd296 : phinc={ 12'd1601 };
        10'd297 : phinc={ 12'd1602 };
        10'd298 : phinc={ 12'd1604 };
        10'd299 : phinc={ 12'd1605 };
        10'd300 : phinc={ 12'd1607 };
        10'd301 : phinc={ 12'd1608 };
        10'd302 : phinc={ 12'd1609 };
        10'd303 : phinc={ 12'd1610 };
        10'd304 : phinc={ 12'd1613 };
        10'd305 : phinc={ 12'd1614 };
        10'd306 : phinc={ 12'd1615 };
        10'd307 : phinc={ 12'd1616 };
        10'd308 : phinc={ 12'd1618 };
        10'd309 : phinc={ 12'd1619 };
        10'd310 : phinc={ 12'd1621 };
        10'd311 : phinc={ 12'd1622 };
        10'd312 : phinc={ 12'd1624 };
        10'd313 : phinc={ 12'd1625 };
        10'd314 : phinc={ 12'd1627 };
        10'd315 : phinc={ 12'd1628 };
        10'd316 : phinc={ 12'd1630 };
        10'd317 : phinc={ 12'd1631 };
        10'd318 : phinc={ 12'd1632 };
        10'd319 : phinc={ 12'd1633 };
        10'd320 : phinc={ 12'd1637 };
        10'd321 : phinc={ 12'd1638 };
        10'd322 : phinc={ 12'd1639 };
        10'd323 : phinc={ 12'd1640 };
        10'd324 : phinc={ 12'd1642 };
        10'd325 : phinc={ 12'd1643 };
        10'd326 : phinc={ 12'd1645 };
        10'd327 : phinc={ 12'd1646 };
        10'd328 : phinc={ 12'd1648 };
        10'd329 : phinc={ 12'd1649 };
        10'd330 : phinc={ 12'd1651 };
        10'd331 : phinc={ 12'd1652 };
        10'd332 : phinc={ 12'd1654 };
        10'd333 : phinc={ 12'd1655 };
        10'd334 : phinc={ 12'd1656 };
        10'd335 : phinc={ 12'd1657 };
        10'd336 : phinc={ 12'd1660 };
        10'd337 : phinc={ 12'd1661 };
        10'd338 : phinc={ 12'd1663 };
        10'd339 : phinc={ 12'd1664 };
        10'd340 : phinc={ 12'd1666 };
        10'd341 : phinc={ 12'd1667 };
        10'd342 : phinc={ 12'd1669 };
        10'd343 : phinc={ 12'd1670 };
        10'd344 : phinc={ 12'd1672 };
        10'd345 : phinc={ 12'd1673 };
        10'd346 : phinc={ 12'd1675 };
        10'd347 : phinc={ 12'd1676 };
        10'd348 : phinc={ 12'd1678 };
        10'd349 : phinc={ 12'd1679 };
        10'd350 : phinc={ 12'd1681 };
        10'd351 : phinc={ 12'd1682 };
        10'd352 : phinc={ 12'd1685 };
        10'd353 : phinc={ 12'd1686 };
        10'd354 : phinc={ 12'd1688 };
        10'd355 : phinc={ 12'd1689 };
        10'd356 : phinc={ 12'd1691 };
        10'd357 : phinc={ 12'd1692 };
        10'd358 : phinc={ 12'd1694 };
        10'd359 : phinc={ 12'd1695 };
        10'd360 : phinc={ 12'd1697 };
        10'd361 : phinc={ 12'd1698 };
        10'd362 : phinc={ 12'd1700 };
        10'd363 : phinc={ 12'd1701 };
        10'd364 : phinc={ 12'd1703 };
        10'd365 : phinc={ 12'd1704 };
        10'd366 : phinc={ 12'd1706 };
        10'd367 : phinc={ 12'd1707 };
        10'd368 : phinc={ 12'd1709 };
        10'd369 : phinc={ 12'd1710 };
        10'd370 : phinc={ 12'd1712 };
        10'd371 : phinc={ 12'd1713 };
        10'd372 : phinc={ 12'd1715 };
        10'd373 : phinc={ 12'd1716 };
        10'd374 : phinc={ 12'd1718 };
        10'd375 : phinc={ 12'd1719 };
        10'd376 : phinc={ 12'd1721 };
        10'd377 : phinc={ 12'd1722 };
        10'd378 : phinc={ 12'd1724 };
        10'd379 : phinc={ 12'd1725 };
        10'd380 : phinc={ 12'd1727 };
        10'd381 : phinc={ 12'd1728 };
        10'd382 : phinc={ 12'd1730 };
        10'd383 : phinc={ 12'd1731 };
        10'd384 : phinc={ 12'd1734 };
        10'd385 : phinc={ 12'd1735 };
        10'd386 : phinc={ 12'd1737 };
        10'd387 : phinc={ 12'd1738 };
        10'd388 : phinc={ 12'd1740 };
        10'd389 : phinc={ 12'd1741 };
        10'd390 : phinc={ 12'd1743 };
        10'd391 : phinc={ 12'd1744 };
        10'd392 : phinc={ 12'd1746 };
        10'd393 : phinc={ 12'd1748 };
        10'd394 : phinc={ 12'd1749 };
        10'd395 : phinc={ 12'd1751 };
        10'd396 : phinc={ 12'd1752 };
        10'd397 : phinc={ 12'd1754 };
        10'd398 : phinc={ 12'd1755 };
        10'd399 : phinc={ 12'd1757 };
        10'd400 : phinc={ 12'd1759 };
        10'd401 : phinc={ 12'd1760 };
        10'd402 : phinc={ 12'd1762 };
        10'd403 : phinc={ 12'd1763 };
        10'd404 : phinc={ 12'd1765 };
        10'd405 : phinc={ 12'd1766 };
        10'd406 : phinc={ 12'd1768 };
        10'd407 : phinc={ 12'd1769 };
        10'd408 : phinc={ 12'd1771 };
        10'd409 : phinc={ 12'd1773 };
        10'd410 : phinc={ 12'd1774 };
        10'd411 : phinc={ 12'd1776 };
        10'd412 : phinc={ 12'd1777 };
        10'd413 : phinc={ 12'd1779 };
        10'd414 : phinc={ 12'd1780 };
        10'd415 : phinc={ 12'd1782 };
        10'd416 : phinc={ 12'd1785 };
        10'd417 : phinc={ 12'd1786 };
        10'd418 : phinc={ 12'd1788 };
        10'd419 : phinc={ 12'd1789 };
        10'd420 : phinc={ 12'd1791 };
        10'd421 : phinc={ 12'd1793 };
        10'd422 : phinc={ 12'd1794 };
        10'd423 : phinc={ 12'd1796 };
        10'd424 : phinc={ 12'd1798 };
        10'd425 : phinc={ 12'd1799 };
        10'd426 : phinc={ 12'd1801 };
        10'd427 : phinc={ 12'd1802 };
        10'd428 : phinc={ 12'd1804 };
        10'd429 : phinc={ 12'd1806 };
        10'd430 : phinc={ 12'd1807 };
        10'd431 : phinc={ 12'd1809 };
        10'd432 : phinc={ 12'd1811 };
        10'd433 : phinc={ 12'd1812 };
        10'd434 : phinc={ 12'd1814 };
        10'd435 : phinc={ 12'd1815 };
        10'd436 : phinc={ 12'd1817 };
        10'd437 : phinc={ 12'd1819 };
        10'd438 : phinc={ 12'd1820 };
        10'd439 : phinc={ 12'd1822 };
        10'd440 : phinc={ 12'd1824 };
        10'd441 : phinc={ 12'd1825 };
        10'd442 : phinc={ 12'd1827 };
        10'd443 : phinc={ 12'd1828 };
        10'd444 : phinc={ 12'd1830 };
        10'd445 : phinc={ 12'd1832 };
        10'd446 : phinc={ 12'd1833 };
        10'd447 : phinc={ 12'd1835 };
        10'd448 : phinc={ 12'd0 };
        10'd449 : phinc={ 12'd2 };
        10'd450 : phinc={ 12'd4 };
        10'd451 : phinc={ 12'd6 };
        10'd452 : phinc={ 12'd4 };
        10'd453 : phinc={ 12'd6 };
        10'd454 : phinc={ 12'd8 };
        10'd455 : phinc={ 12'd10 };
        10'd456 : phinc={ 12'd9 };
        10'd457 : phinc={ 12'd11 };
        10'd458 : phinc={ 12'd13 };
        10'd459 : phinc={ 12'd15 };
        10'd460 : phinc={ 12'd15 };
        10'd461 : phinc={ 12'd17 };
        10'd462 : phinc={ 12'd19 };
        10'd463 : phinc={ 12'd21 };
        10'd464 : phinc={ 12'd0 };
        10'd465 : phinc={ 12'd2 };
        10'd466 : phinc={ 12'd4 };
        10'd467 : phinc={ 12'd6 };
        10'd468 : phinc={ 12'd4 };
        10'd469 : phinc={ 12'd6 };
        10'd470 : phinc={ 12'd8 };
        10'd471 : phinc={ 12'd10 };
        10'd472 : phinc={ 12'd9 };
        10'd473 : phinc={ 12'd11 };
        10'd474 : phinc={ 12'd13 };
        10'd475 : phinc={ 12'd15 };
        10'd476 : phinc={ 12'd15 };
        10'd477 : phinc={ 12'd17 };
        10'd478 : phinc={ 12'd19 };
        10'd479 : phinc={ 12'd21 };
        10'd480 : phinc={ 12'd0 };
        10'd481 : phinc={ 12'd2 };
        10'd482 : phinc={ 12'd4 };
        10'd483 : phinc={ 12'd6 };
        10'd484 : phinc={ 12'd4 };
        10'd485 : phinc={ 12'd6 };
        10'd486 : phinc={ 12'd8 };
        10'd487 : phinc={ 12'd10 };
        10'd488 : phinc={ 12'd9 };
        10'd489 : phinc={ 12'd11 };
        10'd490 : phinc={ 12'd13 };
        10'd491 : phinc={ 12'd15 };
        10'd492 : phinc={ 12'd15 };
        10'd493 : phinc={ 12'd17 };
        10'd494 : phinc={ 12'd19 };
        10'd495 : phinc={ 12'd21 };
        10'd496 : phinc={ 12'd0 };
        10'd497 : phinc={ 12'd2 };
        10'd498 : phinc={ 12'd4 };
        10'd499 : phinc={ 12'd6 };
        10'd500 : phinc={ 12'd4 };
        10'd501 : phinc={ 12'd6 };
        10'd502 : phinc={ 12'd8 };
        10'd503 : phinc={ 12'd10 };
        10'd504 : phinc={ 12'd9 };
        10'd505 : phinc={ 12'd11 };
        10'd506 : phinc={ 12'd13 };
        10'd507 : phinc={ 12'd15 };
        10'd508 : phinc={ 12'd15 };
        10'd509 : phinc={ 12'd17 };
        10'd510 : phinc={ 12'd19 };
        10'd511 : phinc={ 12'd21 };
        10'd512 : phinc={ 12'd1837 };
        10'd513 : phinc={ 12'd1838 };
        10'd514 : phinc={ 12'd1840 };
        10'd515 : phinc={ 12'd1841 };
        10'd516 : phinc={ 12'd1843 };
        10'd517 : phinc={ 12'd1845 };
        10'd518 : phinc={ 12'd1846 };
        10'd519 : phinc={ 12'd1848 };
        10'd520 : phinc={ 12'd1850 };
        10'd521 : phinc={ 12'd1851 };
        10'd522 : phinc={ 12'd1853 };
        10'd523 : phinc={ 12'd1854 };
        10'd524 : phinc={ 12'd1856 };
        10'd525 : phinc={ 12'd1858 };
        10'd526 : phinc={ 12'd1859 };
        10'd527 : phinc={ 12'd1861 };
        10'd528 : phinc={ 12'd1864 };
        10'd529 : phinc={ 12'd1865 };
        10'd530 : phinc={ 12'd1867 };
        10'd531 : phinc={ 12'd1868 };
        10'd532 : phinc={ 12'd1870 };
        10'd533 : phinc={ 12'd1872 };
        10'd534 : phinc={ 12'd1873 };
        10'd535 : phinc={ 12'd1875 };
        10'd536 : phinc={ 12'd1877 };
        10'd537 : phinc={ 12'd1879 };
        10'd538 : phinc={ 12'd1880 };
        10'd539 : phinc={ 12'd1882 };
        10'd540 : phinc={ 12'd1884 };
        10'd541 : phinc={ 12'd1885 };
        10'd542 : phinc={ 12'd1887 };
        10'd543 : phinc={ 12'd1888 };
        10'd544 : phinc={ 12'd1891 };
        10'd545 : phinc={ 12'd1892 };
        10'd546 : phinc={ 12'd1894 };
        10'd547 : phinc={ 12'd1895 };
        10'd548 : phinc={ 12'd1897 };
        10'd549 : phinc={ 12'd1899 };
        10'd550 : phinc={ 12'd1900 };
        10'd551 : phinc={ 12'd1902 };
        10'd552 : phinc={ 12'd1904 };
        10'd553 : phinc={ 12'd1906 };
        10'd554 : phinc={ 12'd1907 };
        10'd555 : phinc={ 12'd1909 };
        10'd556 : phinc={ 12'd1911 };
        10'd557 : phinc={ 12'd1912 };
        10'd558 : phinc={ 12'd1914 };
        10'd559 : phinc={ 12'd1915 };
        10'd560 : phinc={ 12'd1918 };
        10'd561 : phinc={ 12'd1919 };
        10'd562 : phinc={ 12'd1921 };
        10'd563 : phinc={ 12'd1923 };
        10'd564 : phinc={ 12'd1925 };
        10'd565 : phinc={ 12'd1926 };
        10'd566 : phinc={ 12'd1928 };
        10'd567 : phinc={ 12'd1930 };
        10'd568 : phinc={ 12'd1932 };
        10'd569 : phinc={ 12'd1933 };
        10'd570 : phinc={ 12'd1935 };
        10'd571 : phinc={ 12'd1937 };
        10'd572 : phinc={ 12'd1939 };
        10'd573 : phinc={ 12'd1940 };
        10'd574 : phinc={ 12'd1942 };
        10'd575 : phinc={ 12'd1944 };
        10'd576 : phinc={ 12'd1946 };
        10'd577 : phinc={ 12'd1947 };
        10'd578 : phinc={ 12'd1949 };
        10'd579 : phinc={ 12'd1951 };
        10'd580 : phinc={ 12'd1953 };
        10'd581 : phinc={ 12'd1954 };
        10'd582 : phinc={ 12'd1956 };
        10'd583 : phinc={ 12'd1958 };
        10'd584 : phinc={ 12'd1960 };
        10'd585 : phinc={ 12'd1961 };
        10'd586 : phinc={ 12'd1963 };
        10'd587 : phinc={ 12'd1965 };
        10'd588 : phinc={ 12'd1967 };
        10'd589 : phinc={ 12'd1968 };
        10'd590 : phinc={ 12'd1970 };
        10'd591 : phinc={ 12'd1972 };
        10'd592 : phinc={ 12'd1975 };
        10'd593 : phinc={ 12'd1976 };
        10'd594 : phinc={ 12'd1978 };
        10'd595 : phinc={ 12'd1980 };
        10'd596 : phinc={ 12'd1982 };
        10'd597 : phinc={ 12'd1983 };
        10'd598 : phinc={ 12'd1985 };
        10'd599 : phinc={ 12'd1987 };
        10'd600 : phinc={ 12'd1989 };
        10'd601 : phinc={ 12'd1990 };
        10'd602 : phinc={ 12'd1992 };
        10'd603 : phinc={ 12'd1994 };
        10'd604 : phinc={ 12'd1996 };
        10'd605 : phinc={ 12'd1997 };
        10'd606 : phinc={ 12'd1999 };
        10'd607 : phinc={ 12'd2001 };
        10'd608 : phinc={ 12'd2003 };
        10'd609 : phinc={ 12'd2004 };
        10'd610 : phinc={ 12'd2006 };
        10'd611 : phinc={ 12'd2008 };
        10'd612 : phinc={ 12'd2010 };
        10'd613 : phinc={ 12'd2011 };
        10'd614 : phinc={ 12'd2013 };
        10'd615 : phinc={ 12'd2015 };
        10'd616 : phinc={ 12'd2017 };
        10'd617 : phinc={ 12'd2019 };
        10'd618 : phinc={ 12'd2021 };
        10'd619 : phinc={ 12'd2022 };
        10'd620 : phinc={ 12'd2024 };
        10'd621 : phinc={ 12'd2026 };
        10'd622 : phinc={ 12'd2028 };
        10'd623 : phinc={ 12'd2029 };
        10'd624 : phinc={ 12'd2032 };
        10'd625 : phinc={ 12'd2033 };
        10'd626 : phinc={ 12'd2035 };
        10'd627 : phinc={ 12'd2037 };
        10'd628 : phinc={ 12'd2039 };
        10'd629 : phinc={ 12'd2041 };
        10'd630 : phinc={ 12'd2043 };
        10'd631 : phinc={ 12'd2044 };
        10'd632 : phinc={ 12'd2047 };
        10'd633 : phinc={ 12'd2048 };
        10'd634 : phinc={ 12'd2050 };
        10'd635 : phinc={ 12'd2052 };
        10'd636 : phinc={ 12'd2054 };
        10'd637 : phinc={ 12'd2056 };
        10'd638 : phinc={ 12'd2058 };
        10'd639 : phinc={ 12'd2059 };
        10'd640 : phinc={ 12'd2062 };
        10'd641 : phinc={ 12'd2063 };
        10'd642 : phinc={ 12'd2065 };
        10'd643 : phinc={ 12'd2067 };
        10'd644 : phinc={ 12'd2069 };
        10'd645 : phinc={ 12'd2071 };
        10'd646 : phinc={ 12'd2073 };
        10'd647 : phinc={ 12'd2074 };
        10'd648 : phinc={ 12'd2077 };
        10'd649 : phinc={ 12'd2078 };
        10'd650 : phinc={ 12'd2080 };
        10'd651 : phinc={ 12'd2082 };
        10'd652 : phinc={ 12'd2084 };
        10'd653 : phinc={ 12'd2086 };
        10'd654 : phinc={ 12'd2088 };
        10'd655 : phinc={ 12'd2089 };
        10'd656 : phinc={ 12'd2092 };
        10'd657 : phinc={ 12'd2093 };
        10'd658 : phinc={ 12'd2095 };
        10'd659 : phinc={ 12'd2097 };
        10'd660 : phinc={ 12'd2099 };
        10'd661 : phinc={ 12'd2101 };
        10'd662 : phinc={ 12'd2103 };
        10'd663 : phinc={ 12'd2104 };
        10'd664 : phinc={ 12'd2107 };
        10'd665 : phinc={ 12'd2108 };
        10'd666 : phinc={ 12'd2110 };
        10'd667 : phinc={ 12'd2112 };
        10'd668 : phinc={ 12'd2114 };
        10'd669 : phinc={ 12'd2116 };
        10'd670 : phinc={ 12'd2118 };
        10'd671 : phinc={ 12'd2119 };
        10'd672 : phinc={ 12'd2122 };
        10'd673 : phinc={ 12'd2123 };
        10'd674 : phinc={ 12'd2125 };
        10'd675 : phinc={ 12'd2127 };
        10'd676 : phinc={ 12'd2129 };
        10'd677 : phinc={ 12'd2131 };
        10'd678 : phinc={ 12'd2133 };
        10'd679 : phinc={ 12'd2134 };
        10'd680 : phinc={ 12'd2137 };
        10'd681 : phinc={ 12'd2139 };
        10'd682 : phinc={ 12'd2141 };
        10'd683 : phinc={ 12'd2142 };
        10'd684 : phinc={ 12'd2145 };
        10'd685 : phinc={ 12'd2146 };
        10'd686 : phinc={ 12'd2148 };
        10'd687 : phinc={ 12'd2150 };
        10'd688 : phinc={ 12'd2153 };
        10'd689 : phinc={ 12'd2154 };
        10'd690 : phinc={ 12'd2156 };
        10'd691 : phinc={ 12'd2158 };
        10'd692 : phinc={ 12'd2160 };
        10'd693 : phinc={ 12'd2162 };
        10'd694 : phinc={ 12'd2164 };
        10'd695 : phinc={ 12'd2165 };
        10'd696 : phinc={ 12'd2168 };
        10'd697 : phinc={ 12'd2170 };
        10'd698 : phinc={ 12'd2172 };
        10'd699 : phinc={ 12'd2173 };
        10'd700 : phinc={ 12'd2176 };
        10'd701 : phinc={ 12'd2177 };
        10'd702 : phinc={ 12'd2179 };
        10'd703 : phinc={ 12'd2181 };
        10'd704 : phinc={ 12'd0 };
        10'd705 : phinc={ 12'd2 };
        10'd706 : phinc={ 12'd4 };
        10'd707 : phinc={ 12'd6 };
        10'd708 : phinc={ 12'd4 };
        10'd709 : phinc={ 12'd6 };
        10'd710 : phinc={ 12'd8 };
        10'd711 : phinc={ 12'd10 };
        10'd712 : phinc={ 12'd9 };
        10'd713 : phinc={ 12'd11 };
        10'd714 : phinc={ 12'd13 };
        10'd715 : phinc={ 12'd15 };
        10'd716 : phinc={ 12'd15 };
        10'd717 : phinc={ 12'd17 };
        10'd718 : phinc={ 12'd19 };
        10'd719 : phinc={ 12'd21 };
        10'd720 : phinc={ 12'd0 };
        10'd721 : phinc={ 12'd2 };
        10'd722 : phinc={ 12'd4 };
        10'd723 : phinc={ 12'd6 };
        10'd724 : phinc={ 12'd4 };
        10'd725 : phinc={ 12'd6 };
        10'd726 : phinc={ 12'd8 };
        10'd727 : phinc={ 12'd10 };
        10'd728 : phinc={ 12'd9 };
        10'd729 : phinc={ 12'd11 };
        10'd730 : phinc={ 12'd13 };
        10'd731 : phinc={ 12'd15 };
        10'd732 : phinc={ 12'd15 };
        10'd733 : phinc={ 12'd17 };
        10'd734 : phinc={ 12'd19 };
        10'd735 : phinc={ 12'd21 };
        10'd736 : phinc={ 12'd0 };
        10'd737 : phinc={ 12'd2 };
        10'd738 : phinc={ 12'd4 };
        10'd739 : phinc={ 12'd6 };
        10'd740 : phinc={ 12'd4 };
        10'd741 : phinc={ 12'd6 };
        10'd742 : phinc={ 12'd8 };
        10'd743 : phinc={ 12'd10 };
        10'd744 : phinc={ 12'd9 };
        10'd745 : phinc={ 12'd11 };
        10'd746 : phinc={ 12'd13 };
        10'd747 : phinc={ 12'd15 };
        10'd748 : phinc={ 12'd15 };
        10'd749 : phinc={ 12'd17 };
        10'd750 : phinc={ 12'd19 };
        10'd751 : phinc={ 12'd21 };
        10'd752 : phinc={ 12'd0 };
        10'd753 : phinc={ 12'd2 };
        10'd754 : phinc={ 12'd4 };
        10'd755 : phinc={ 12'd6 };
        10'd756 : phinc={ 12'd4 };
        10'd757 : phinc={ 12'd6 };
        10'd758 : phinc={ 12'd8 };
        10'd759 : phinc={ 12'd10 };
        10'd760 : phinc={ 12'd9 };
        10'd761 : phinc={ 12'd11 };
        10'd762 : phinc={ 12'd13 };
        10'd763 : phinc={ 12'd15 };
        10'd764 : phinc={ 12'd15 };
        10'd765 : phinc={ 12'd17 };
        10'd766 : phinc={ 12'd19 };
        10'd767 : phinc={ 12'd21 };
        10'd768 : phinc={ 12'd2185 };
        10'd769 : phinc={ 12'd2186 };
        10'd770 : phinc={ 12'd2188 };
        10'd771 : phinc={ 12'd2190 };
        10'd772 : phinc={ 12'd2192 };
        10'd773 : phinc={ 12'd2194 };
        10'd774 : phinc={ 12'd2196 };
        10'd775 : phinc={ 12'd2197 };
        10'd776 : phinc={ 12'd2200 };
        10'd777 : phinc={ 12'd2202 };
        10'd778 : phinc={ 12'd2204 };
        10'd779 : phinc={ 12'd2205 };
        10'd780 : phinc={ 12'd2208 };
        10'd781 : phinc={ 12'd2209 };
        10'd782 : phinc={ 12'd2211 };
        10'd783 : phinc={ 12'd2213 };
        10'd784 : phinc={ 12'd2216 };
        10'd785 : phinc={ 12'd2218 };
        10'd786 : phinc={ 12'd2220 };
        10'd787 : phinc={ 12'd2222 };
        10'd788 : phinc={ 12'd2223 };
        10'd789 : phinc={ 12'd2226 };
        10'd790 : phinc={ 12'd2227 };
        10'd791 : phinc={ 12'd2230 };
        10'd792 : phinc={ 12'd2232 };
        10'd793 : phinc={ 12'd2234 };
        10'd794 : phinc={ 12'd2236 };
        10'd795 : phinc={ 12'd2238 };
        10'd796 : phinc={ 12'd2239 };
        10'd797 : phinc={ 12'd2242 };
        10'd798 : phinc={ 12'd2243 };
        10'd799 : phinc={ 12'd2246 };
        10'd800 : phinc={ 12'd2249 };
        10'd801 : phinc={ 12'd2251 };
        10'd802 : phinc={ 12'd2253 };
        10'd803 : phinc={ 12'd2255 };
        10'd804 : phinc={ 12'd2256 };
        10'd805 : phinc={ 12'd2259 };
        10'd806 : phinc={ 12'd2260 };
        10'd807 : phinc={ 12'd2263 };
        10'd808 : phinc={ 12'd2265 };
        10'd809 : phinc={ 12'd2267 };
        10'd810 : phinc={ 12'd2269 };
        10'd811 : phinc={ 12'd2271 };
        10'd812 : phinc={ 12'd2272 };
        10'd813 : phinc={ 12'd2275 };
        10'd814 : phinc={ 12'd2276 };
        10'd815 : phinc={ 12'd2279 };
        10'd816 : phinc={ 12'd2281 };
        10'd817 : phinc={ 12'd2283 };
        10'd818 : phinc={ 12'd2285 };
        10'd819 : phinc={ 12'd2287 };
        10'd820 : phinc={ 12'd2288 };
        10'd821 : phinc={ 12'd2291 };
        10'd822 : phinc={ 12'd2292 };
        10'd823 : phinc={ 12'd2295 };
        10'd824 : phinc={ 12'd2297 };
        10'd825 : phinc={ 12'd2299 };
        10'd826 : phinc={ 12'd2301 };
        10'd827 : phinc={ 12'd2303 };
        10'd828 : phinc={ 12'd2304 };
        10'd829 : phinc={ 12'd2307 };
        10'd830 : phinc={ 12'd2308 };
        10'd831 : phinc={ 12'd2311 };
        10'd832 : phinc={ 12'd2315 };
        10'd833 : phinc={ 12'd2317 };
        10'd834 : phinc={ 12'd2319 };
        10'd835 : phinc={ 12'd2321 };
        10'd836 : phinc={ 12'd2322 };
        10'd837 : phinc={ 12'd2325 };
        10'd838 : phinc={ 12'd2326 };
        10'd839 : phinc={ 12'd2329 };
        10'd840 : phinc={ 12'd2331 };
        10'd841 : phinc={ 12'd2333 };
        10'd842 : phinc={ 12'd2335 };
        10'd843 : phinc={ 12'd2337 };
        10'd844 : phinc={ 12'd2338 };
        10'd845 : phinc={ 12'd2341 };
        10'd846 : phinc={ 12'd2342 };
        10'd847 : phinc={ 12'd2345 };
        10'd848 : phinc={ 12'd2348 };
        10'd849 : phinc={ 12'd2350 };
        10'd850 : phinc={ 12'd2352 };
        10'd851 : phinc={ 12'd2354 };
        10'd852 : phinc={ 12'd2355 };
        10'd853 : phinc={ 12'd2358 };
        10'd854 : phinc={ 12'd2359 };
        10'd855 : phinc={ 12'd2362 };
        10'd856 : phinc={ 12'd2364 };
        10'd857 : phinc={ 12'd2366 };
        10'd858 : phinc={ 12'd2368 };
        10'd859 : phinc={ 12'd2370 };
        10'd860 : phinc={ 12'd2371 };
        10'd861 : phinc={ 12'd2374 };
        10'd862 : phinc={ 12'd2375 };
        10'd863 : phinc={ 12'd2378 };
        10'd864 : phinc={ 12'd2382 };
        10'd865 : phinc={ 12'd2384 };
        10'd866 : phinc={ 12'd2386 };
        10'd867 : phinc={ 12'd2388 };
        10'd868 : phinc={ 12'd2389 };
        10'd869 : phinc={ 12'd2392 };
        10'd870 : phinc={ 12'd2393 };
        10'd871 : phinc={ 12'd2396 };
        10'd872 : phinc={ 12'd2398 };
        10'd873 : phinc={ 12'd2400 };
        10'd874 : phinc={ 12'd2402 };
        10'd875 : phinc={ 12'd2404 };
        10'd876 : phinc={ 12'd2407 };
        10'd877 : phinc={ 12'd2410 };
        10'd878 : phinc={ 12'd2411 };
        10'd879 : phinc={ 12'd2414 };
        10'd880 : phinc={ 12'd2417 };
        10'd881 : phinc={ 12'd2419 };
        10'd882 : phinc={ 12'd2421 };
        10'd883 : phinc={ 12'd2423 };
        10'd884 : phinc={ 12'd2424 };
        10'd885 : phinc={ 12'd2427 };
        10'd886 : phinc={ 12'd2428 };
        10'd887 : phinc={ 12'd2431 };
        10'd888 : phinc={ 12'd2433 };
        10'd889 : phinc={ 12'd2435 };
        10'd890 : phinc={ 12'd2437 };
        10'd891 : phinc={ 12'd2439 };
        10'd892 : phinc={ 12'd2442 };
        10'd893 : phinc={ 12'd2445 };
        10'd894 : phinc={ 12'd2446 };
        10'd895 : phinc={ 12'd2449 };
        10'd896 : phinc={ 12'd2452 };
        10'd897 : phinc={ 12'd2454 };
        10'd898 : phinc={ 12'd2456 };
        10'd899 : phinc={ 12'd2458 };
        10'd900 : phinc={ 12'd2459 };
        10'd901 : phinc={ 12'd2462 };
        10'd902 : phinc={ 12'd2463 };
        10'd903 : phinc={ 12'd2466 };
        10'd904 : phinc={ 12'd2468 };
        10'd905 : phinc={ 12'd2470 };
        10'd906 : phinc={ 12'd2472 };
        10'd907 : phinc={ 12'd2474 };
        10'd908 : phinc={ 12'd2477 };
        10'd909 : phinc={ 12'd2480 };
        10'd910 : phinc={ 12'd2481 };
        10'd911 : phinc={ 12'd2484 };
        10'd912 : phinc={ 12'd2488 };
        10'd913 : phinc={ 12'd2490 };
        10'd914 : phinc={ 12'd2492 };
        10'd915 : phinc={ 12'd2494 };
        10'd916 : phinc={ 12'd2495 };
        10'd917 : phinc={ 12'd2498 };
        10'd918 : phinc={ 12'd2499 };
        10'd919 : phinc={ 12'd2502 };
        10'd920 : phinc={ 12'd2504 };
        10'd921 : phinc={ 12'd2506 };
        10'd922 : phinc={ 12'd2508 };
        10'd923 : phinc={ 12'd2510 };
        10'd924 : phinc={ 12'd2513 };
        10'd925 : phinc={ 12'd2516 };
        10'd926 : phinc={ 12'd2517 };
        10'd927 : phinc={ 12'd2520 };
        10'd928 : phinc={ 12'd2524 };
        10'd929 : phinc={ 12'd2526 };
        10'd930 : phinc={ 12'd2528 };
        10'd931 : phinc={ 12'd2530 };
        10'd932 : phinc={ 12'd2531 };
        10'd933 : phinc={ 12'd2534 };
        10'd934 : phinc={ 12'd2535 };
        10'd935 : phinc={ 12'd2538 };
        10'd936 : phinc={ 12'd2540 };
        10'd937 : phinc={ 12'd2542 };
        10'd938 : phinc={ 12'd2544 };
        10'd939 : phinc={ 12'd2546 };
        10'd940 : phinc={ 12'd2549 };
        10'd941 : phinc={ 12'd2552 };
        10'd942 : phinc={ 12'd2553 };
        10'd943 : phinc={ 12'd2556 };
        10'd944 : phinc={ 12'd2561 };
        10'd945 : phinc={ 12'd2563 };
        10'd946 : phinc={ 12'd2565 };
        10'd947 : phinc={ 12'd2567 };
        10'd948 : phinc={ 12'd2568 };
        10'd949 : phinc={ 12'd2571 };
        10'd950 : phinc={ 12'd2572 };
        10'd951 : phinc={ 12'd2575 };
        10'd952 : phinc={ 12'd2577 };
        10'd953 : phinc={ 12'd2579 };
        10'd954 : phinc={ 12'd2581 };
        10'd955 : phinc={ 12'd2583 };
        10'd956 : phinc={ 12'd2586 };
        10'd957 : phinc={ 12'd2589 };
        10'd958 : phinc={ 12'd2590 };
        10'd959 : phinc={ 12'd2593 };
        10'd960 : phinc={ 12'd0 };
        10'd961 : phinc={ 12'd2 };
        10'd962 : phinc={ 12'd4 };
        10'd963 : phinc={ 12'd6 };
        10'd964 : phinc={ 12'd4 };
        10'd965 : phinc={ 12'd6 };
        10'd966 : phinc={ 12'd8 };
        10'd967 : phinc={ 12'd10 };
        10'd968 : phinc={ 12'd9 };
        10'd969 : phinc={ 12'd11 };
        10'd970 : phinc={ 12'd13 };
        10'd971 : phinc={ 12'd15 };
        10'd972 : phinc={ 12'd15 };
        10'd973 : phinc={ 12'd17 };
        10'd974 : phinc={ 12'd19 };
        10'd975 : phinc={ 12'd21 };
        10'd976 : phinc={ 12'd0 };
        10'd977 : phinc={ 12'd2 };
        10'd978 : phinc={ 12'd4 };
        10'd979 : phinc={ 12'd6 };
        10'd980 : phinc={ 12'd4 };
        10'd981 : phinc={ 12'd6 };
        10'd982 : phinc={ 12'd8 };
        10'd983 : phinc={ 12'd10 };
        10'd984 : phinc={ 12'd9 };
        10'd985 : phinc={ 12'd11 };
        10'd986 : phinc={ 12'd13 };
        10'd987 : phinc={ 12'd15 };
        10'd988 : phinc={ 12'd15 };
        10'd989 : phinc={ 12'd17 };
        10'd990 : phinc={ 12'd19 };
        10'd991 : phinc={ 12'd21 };
        10'd992 : phinc={ 12'd0 };
        10'd993 : phinc={ 12'd2 };
        10'd994 : phinc={ 12'd4 };
        10'd995 : phinc={ 12'd6 };
        10'd996 : phinc={ 12'd4 };
        10'd997 : phinc={ 12'd6 };
        10'd998 : phinc={ 12'd8 };
        10'd999 : phinc={ 12'd10 };
        10'd1000: phinc={ 12'd9 };
        10'd1001: phinc={ 12'd11 };
        10'd1002: phinc={ 12'd13 };
        10'd1003: phinc={ 12'd15 };
        10'd1004: phinc={ 12'd15 };
        10'd1005: phinc={ 12'd17 };
        10'd1006: phinc={ 12'd19 };
        10'd1007: phinc={ 12'd21 };
        10'd1008: phinc={ 12'd0 };
        10'd1009: phinc={ 12'd2 };
        10'd1010: phinc={ 12'd4 };
        10'd1011: phinc={ 12'd6 };
        10'd1012: phinc={ 12'd4 };
        10'd1013: phinc={ 12'd6 };
        10'd1014: phinc={ 12'd8 };
        10'd1015: phinc={ 12'd10 };
        10'd1016: phinc={ 12'd9 };
        10'd1017: phinc={ 12'd11 };
        10'd1018: phinc={ 12'd13 };
        10'd1019: phinc={ 12'd15 };
        10'd1020: phinc={ 12'd15 };
        10'd1021: phinc={ 12'd17 };
        10'd1022: phinc={ 12'd19 };
        10'd1023: phinc={ 12'd21 };
    endcase
end

endmodule
